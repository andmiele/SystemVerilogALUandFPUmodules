//-----------------------------------------------------------------------------
// Copyright 2021 Andrea Miele
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------------------

// halfAdder.sv
// sum = x ^ y = (x | y) & (!(x & y)); x,y -> sum: 5 gate-delays
// cout = (x & y); x,y -> cout: 2 gate-delays

module halfAdder
(
    input logic x,
    input logic y,
    output logic sum,
    output logic cout
);

assign sum = x ^ y;
assign cout = (x & y);
endmodule
