//-----------------------------------------------------------------------------
// Copyright 2021 Andrea Miele
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------------------

// Radix4PLA1.sv
// PLA for 1-st quotient bit selection 

module Radix4PLA1
(
input logic [5 : 0] r6Abs,
input logic [3 : 0] y4,
output logic q1
);

always_comb
begin

case ({r6Abs, y4})
10'b0011010000: q1 = 1'b1;
10'b0011100000: q1 = 1'b1;
10'b0011110000: q1 = 1'b1;
10'b0100000000: q1 = 1'b1;
10'b0100010000: q1 = 1'b1;
10'b0100100000: q1 = 1'b1;
10'b0100110000: q1 = 1'b1;
10'b0101000000: q1 = 1'b1;
10'b0101010000: q1 = 1'b1;
10'b0101100000: q1 = 1'b1;
10'b0011100001: q1 = 1'b1;
10'b0011110001: q1 = 1'b1;
10'b0100000001: q1 = 1'b1;
10'b0100010001: q1 = 1'b1;
10'b0100100001: q1 = 1'b1;
10'b0100110001: q1 = 1'b1;
10'b0101000001: q1 = 1'b1;
10'b0101010001: q1 = 1'b1;
10'b0101100001: q1 = 1'b1;
10'b0101110001: q1 = 1'b1;
10'b0011110010: q1 = 1'b1;
10'b0100000010: q1 = 1'b1;
10'b0100010010: q1 = 1'b1;
10'b0100100010: q1 = 1'b1;
10'b0100110010: q1 = 1'b1;
10'b0101000010: q1 = 1'b1;
10'b0101010010: q1 = 1'b1;
10'b0101100010: q1 = 1'b1;
10'b0101110010: q1 = 1'b1;
10'b0110000010: q1 = 1'b1;
10'b0011110011: q1 = 1'b1;
10'b0100000011: q1 = 1'b1;
10'b0100010011: q1 = 1'b1;
10'b0100100011: q1 = 1'b1;
10'b0100110011: q1 = 1'b1;
10'b0101000011: q1 = 1'b1;
10'b0101010011: q1 = 1'b1;
10'b0101100011: q1 = 1'b1;
10'b0101110011: q1 = 1'b1;
10'b0110000011: q1 = 1'b1;
10'b0110010011: q1 = 1'b1;
10'b0110100011: q1 = 1'b1;
10'b0100000100: q1 = 1'b1;
10'b0100010100: q1 = 1'b1;
10'b0100100100: q1 = 1'b1;
10'b0100110100: q1 = 1'b1;
10'b0101000100: q1 = 1'b1;
10'b0101010100: q1 = 1'b1;
10'b0101100100: q1 = 1'b1;
10'b0101110100: q1 = 1'b1;
10'b0110000100: q1 = 1'b1;
10'b0110010100: q1 = 1'b1;
10'b0110100100: q1 = 1'b1;
10'b0110110100: q1 = 1'b1;
10'b0100010101: q1 = 1'b1;
10'b0100100101: q1 = 1'b1;
10'b0100110101: q1 = 1'b1;
10'b0101000101: q1 = 1'b1;
10'b0101010101: q1 = 1'b1;
10'b0101100101: q1 = 1'b1;
10'b0101110101: q1 = 1'b1;
10'b0110000101: q1 = 1'b1;
10'b0110010101: q1 = 1'b1;
10'b0110100101: q1 = 1'b1;
10'b0110110101: q1 = 1'b1;
10'b0111000101: q1 = 1'b1;
10'b0111010101: q1 = 1'b1;
10'b0100100110: q1 = 1'b1;
10'b0100110110: q1 = 1'b1;
10'b0101000110: q1 = 1'b1;
10'b0101010110: q1 = 1'b1;
10'b0101100110: q1 = 1'b1;
10'b0101110110: q1 = 1'b1;
10'b0110000110: q1 = 1'b1;
10'b0110010110: q1 = 1'b1;
10'b0110100110: q1 = 1'b1;
10'b0110110110: q1 = 1'b1;
10'b0111000110: q1 = 1'b1;
10'b0111010110: q1 = 1'b1;
10'b0111100110: q1 = 1'b1;
10'b0100110111: q1 = 1'b1;
10'b0101000111: q1 = 1'b1;
10'b0101010111: q1 = 1'b1;
10'b0101100111: q1 = 1'b1;
10'b0101110111: q1 = 1'b1;
10'b0110000111: q1 = 1'b1;
10'b0110010111: q1 = 1'b1;
10'b0110100111: q1 = 1'b1;
10'b0110110111: q1 = 1'b1;
10'b0111000111: q1 = 1'b1;
10'b0111010111: q1 = 1'b1;
10'b0111100111: q1 = 1'b1;
10'b0111110111: q1 = 1'b1;
10'b0101001000: q1 = 1'b1;
10'b0101011000: q1 = 1'b1;
10'b0101101000: q1 = 1'b1;
10'b0101111000: q1 = 1'b1;
10'b0110001000: q1 = 1'b1;
10'b0110011000: q1 = 1'b1;
10'b0110101000: q1 = 1'b1;
10'b0110111000: q1 = 1'b1;
10'b0111001000: q1 = 1'b1;
10'b0111011000: q1 = 1'b1;
10'b0111101000: q1 = 1'b1;
10'b0111111000: q1 = 1'b1;
10'b1000001000: q1 = 1'b1;
10'b1000011000: q1 = 1'b1;
10'b0101011001: q1 = 1'b1;
10'b0101101001: q1 = 1'b1;
10'b0101111001: q1 = 1'b1;
10'b0110001001: q1 = 1'b1;
10'b0110011001: q1 = 1'b1;
10'b0110101001: q1 = 1'b1;
10'b0110111001: q1 = 1'b1;
10'b0111001001: q1 = 1'b1;
10'b0111011001: q1 = 1'b1;
10'b0111101001: q1 = 1'b1;
10'b0111111001: q1 = 1'b1;
10'b1000001001: q1 = 1'b1;
10'b1000011001: q1 = 1'b1;
10'b1000101001: q1 = 1'b1;
10'b0101011010: q1 = 1'b1;
10'b0101101010: q1 = 1'b1;
10'b0101111010: q1 = 1'b1;
10'b0110001010: q1 = 1'b1;
10'b0110011010: q1 = 1'b1;
10'b0110101010: q1 = 1'b1;
10'b0110111010: q1 = 1'b1;
10'b0111001010: q1 = 1'b1;
10'b0111011010: q1 = 1'b1;
10'b0111101010: q1 = 1'b1;
10'b0111111010: q1 = 1'b1;
10'b1000001010: q1 = 1'b1;
10'b1000011010: q1 = 1'b1;
10'b1000101010: q1 = 1'b1;
10'b1000111010: q1 = 1'b1;
10'b0101101011: q1 = 1'b1;
10'b0101111011: q1 = 1'b1;
10'b0110001011: q1 = 1'b1;
10'b0110011011: q1 = 1'b1;
10'b0110101011: q1 = 1'b1;
10'b0110111011: q1 = 1'b1;
10'b0111001011: q1 = 1'b1;
10'b0111011011: q1 = 1'b1;
10'b0111101011: q1 = 1'b1;
10'b0111111011: q1 = 1'b1;
10'b1000001011: q1 = 1'b1;
10'b1000011011: q1 = 1'b1;
10'b1000101011: q1 = 1'b1;
10'b1000111011: q1 = 1'b1;
10'b1001001011: q1 = 1'b1;
10'b1001011011: q1 = 1'b1;
10'b0101111100: q1 = 1'b1;
10'b0110001100: q1 = 1'b1;
10'b0110011100: q1 = 1'b1;
10'b0110101100: q1 = 1'b1;
10'b0110111100: q1 = 1'b1;
10'b0111001100: q1 = 1'b1;
10'b0111011100: q1 = 1'b1;
10'b0111101100: q1 = 1'b1;
10'b0111111100: q1 = 1'b1;
10'b1000001100: q1 = 1'b1;
10'b1000011100: q1 = 1'b1;
10'b1000101100: q1 = 1'b1;
10'b1000111100: q1 = 1'b1;
10'b1001001100: q1 = 1'b1;
10'b1001011100: q1 = 1'b1;
10'b1001101100: q1 = 1'b1;
10'b0110001101: q1 = 1'b1;
10'b0110011101: q1 = 1'b1;
10'b0110101101: q1 = 1'b1;
10'b0110111101: q1 = 1'b1;
10'b0111001101: q1 = 1'b1;
10'b0111011101: q1 = 1'b1;
10'b0111101101: q1 = 1'b1;
10'b0111111101: q1 = 1'b1;
10'b1000001101: q1 = 1'b1;
10'b1000011101: q1 = 1'b1;
10'b1000101101: q1 = 1'b1;
10'b1000111101: q1 = 1'b1;
10'b1001001101: q1 = 1'b1;
10'b1001011101: q1 = 1'b1;
10'b1001101101: q1 = 1'b1;
10'b1001111101: q1 = 1'b1;
10'b0110001110: q1 = 1'b1;
10'b0110011110: q1 = 1'b1;
10'b0110101110: q1 = 1'b1;
10'b0110111110: q1 = 1'b1;
10'b0111001110: q1 = 1'b1;
10'b0111011110: q1 = 1'b1;
10'b0111101110: q1 = 1'b1;
10'b0111111110: q1 = 1'b1;
10'b1000001110: q1 = 1'b1;
10'b1000011110: q1 = 1'b1;
10'b1000101110: q1 = 1'b1;
10'b1000111110: q1 = 1'b1;
10'b1001001110: q1 = 1'b1;
10'b1001011110: q1 = 1'b1;
10'b1001101110: q1 = 1'b1;
10'b1001111110: q1 = 1'b1;
10'b1010001110: q1 = 1'b1;
10'b1010011110: q1 = 1'b1;
10'b0110011111: q1 = 1'b1;
10'b0110101111: q1 = 1'b1;
10'b0110111111: q1 = 1'b1;
10'b0111001111: q1 = 1'b1;
10'b0111011111: q1 = 1'b1;
10'b0111101111: q1 = 1'b1;
10'b0111111111: q1 = 1'b1;
10'b1000001111: q1 = 1'b1;
10'b1000011111: q1 = 1'b1;
10'b1000101111: q1 = 1'b1;
10'b1000111111: q1 = 1'b1;
10'b1001001111: q1 = 1'b1;
10'b1001011111: q1 = 1'b1;
10'b1001101111: q1 = 1'b1;
10'b1001111111: q1 = 1'b1;
10'b1010001111: q1 = 1'b1;
10'b1010011111: q1 = 1'b1;
10'b1010101111: q1 = 1'b1;
default:        q1 = 1'b0;
endcase
end

endmodule
