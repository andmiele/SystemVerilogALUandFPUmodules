//-----------------------------------------------------------------------------
// Copyright 2022 Andrea Miele
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
//-----------------------------------------------------------------------------

// prefixAddSub.sv
// prefix/scan Adder-Subtractor

// Addition with carry propagation computed as parallel prefix-tree for carry propagate (p)
// and generate(p) signals.
// Each node of the prefix-tree is either a pass-through: p_out = p_in and g_out = g_in
// or an operator node: p_out = p1 & p2, g_out = (g1 & p2) | g2
// The critical path for an M-bit adder is about 2 * log_2(M) nodes and the number of gates is
// O(M * log_2(M))
// At level 0 of the tree g and p signals are generated by the M full-adders adding the input bits.
// There are an up-sweep phase and a down-sweep phase.
// In the up-sweep phase there are ceiling(log_2(M)) and at level i (for i = 1 to ceiling(log_2(M))) the previous level horizontal indices of the input pairs
// (p1,p2) and (g1, g2) to the operator nodes are (j * 2**i - 2**(i - 1) - 1, j * 2**i - 1) with the left index being also
// the output index (for all the other indices a pass-through node is used)
// In the down-sweep phase there are ceiling(log_2(M)) - 1 levels and at level i (ceiling(log_2(M)) - 1 down to 1)
// the horizontal indices of the input pairs
// (p1,p2) and (g1, g2) to the operator nodes are (j * 2**i + 2**(i - 1) - 1, j * 2**i - 1) with the left index being also
// the output index (for all the other indices a pass-through node is used)
// See https://en.wikipedia.org/wiki/Prefix_sum for more info on parallel prefix-tree computations 


// Each node of the tree 

module pgOp
(
    input logic g1,
    input logic p1,
    input logic g2,
    input logic p2,
    output logic g,
    output logic p
);
assign g = (g1 & p2) | g2;
assign p = p1 & p2;
endmodule

module fullAdderPGC
(
    input logic cin,
    input logic x,
    input logic y,
    output logic sum,
    output logic g,
    output logic p
);
assign p = x ^ y;
assign g = x & y;
assign sum = p ^ cin;

endmodule

module prefixAddSub
#(parameter M = 32)
(
    input logic sub,
    input logic cin, // arithmetic carry ignored if sub is 1
    input logic [M - 1 : 0] x,
    input logic [M - 1 : 0] y,
    output logic [M - 1 : 0] out,
    output logic cout,
    output logic v
);

localparam N_LVLS = $clog2(M);

logic [M - 1 : 0] yn;
logic [M - 1 : 0] sumi;
logic [M - 1 : 0] p_up [0 : N_LVLS];
logic [M - 1 : 0] g_up [0 : N_LVLS];
logic [M - 1 : 0] p_down [1 : N_LVLS];
logic [M - 1 : 0] g_down [1 : N_LVLS];

logic g0, p0;
assign yn = y ^ {(M){sub}};

assign g_down[N_LVLS] = g_up[N_LVLS];
assign p_down[N_LVLS] = p_up[N_LVLS];

// level 0

// FA0
fullAdderPGC fa_0_0(.cin(sub | cin), .x(x[0]), .y(yn[0]),
    .sum(sumi[0]), .g(g0), 
.p(p0));

assign g_up[0][0] = g0 | (p0 & (sub | cin));
assign p_up[0][0] = 1'b1;

genvar i, j;
generate
for(i = 1; i < M; i++)
begin: lv_0
    fullAdderPGC fa_0_i(.cin(1'b0), .x(x[i]), .y(yn[i]),
        .sum(sumi[i]), .g(g_up[0][i]), 
    .p(p_up[0][i]));
end


// UP-SWEEP
// levels 1 - N_LVLS

for(i = 1; i <= N_LVLS; i++)
begin: lv_i_up
    for(j = 2**i; j <= M; j = j + 2**i)
    begin: lv_j_up
        pgOp op_i_j_up(
            .g1(g_up[i - 1][j - 1 - 2**(i - 1)]), 
            .p1(p_up[i - 1][j - 1 - 2**(i - 1)]),
            .g2(g_up[i - 1][j - 1]), 
            .p2(p_up[i - 1][j - 1]),
            .g(g_up[i][j - 1]), 
        .p(p_up[i][j - 1]));
    end

    // pass-through, j not divisible by 2**I or equal to 0
    for(j = 0; j < M; j = j + 1)
    begin: lv_i_pass_up
        if (((j + 1) % (2**i)) | (j == 0))
        begin: pass_up_if   
            assign g_up[i][j] = g_up[i - 1][j];
            assign p_up[i][j] = p_up[i - 1][j];
        end
    end

end

// DOWN-SWEEP
// levels (N_LVLS - 1) - 1

for(i = N_LVLS - 1; i > 0; i--)
begin: lv_i_down
    for(j = 2**i; j < M - 2**(i - 1); j = j + 2**i)
    begin: lv_j_down   
        pgOp op_i_j_down(
            .g1(g_down[i + 1][j - 1]), 
            .p1(p_down[i + 1][j - 1]),
            .g2(g_down[i + 1][j - 1 + 2**(i - 1)]), 
            .p2(p_down[i + 1][j - 1 + 2**(i - 1)]),
            .g(g_down[i][j - 1 + 2**(i - 1)]), 
        .p(p_down[i][j - 1 + 2**(i - 1)]));
    end

    // pass-through
    for(j = 0; j < M; j = j + 1)
    begin: lv_i_pass_down
        if (!((j >= 2**i) && (j % 2**i == (2**i + 2**(i-1) - 1) % 2**i)))
        begin: pass_down_if   
            assign g_down[i][j] = g_down[i + 1][j];
            assign p_down[i][j] = p_down[i + 1][j];
        end
    end

end
endgenerate

assign cout = g_down[1][M - 1];
assign v = g_down[1][M - 1] ^ g_down[1][M - 2];

assign out[0] = sumi[0];
assign out[M - 1 : 1] = sumi[M - 1 : 1] ^ g_down[1][M - 2 : 0];

endmodule
